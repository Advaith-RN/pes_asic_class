module mult8 (input [2:0] a, output [5:0] y);
	assign y = a*9;
endmodule
